
module Simple (
  // input
  input clk,
  input rst_n
);

endmodule
